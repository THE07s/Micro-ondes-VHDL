library ieee;
use ieee.std_logic_1164.all;

entity micro-ondes is
  port(
    port(
      clk_i, reset_i : in std_logic;
      
  )
