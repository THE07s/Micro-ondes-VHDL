library ieee;
use ieee.std_logic_1164.all;

entity micro-ondes is
  port(
    port        : in std_logic;
  )
